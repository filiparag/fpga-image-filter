package CustomTypes is

    constant kernel_dimension    : integer := 15;
    constant image_slice_width   : integer := 256;
    constant image_slice_height  : integer := 15;

    type flag			    is STD_LOGIC;
    type pixel 		        is array (7 downto 0) 					        of STD_LOGIC;
    type image_slice_row    is array ((image_slice_width - 1) downto 0)     of pixel;
    type kernel_slice_row   is array ((kernel_dimension - 1) downto 0) 	    of pixel;
    type image_slice	    is array ((image_slice_height - 1) downto 0)    of image_slice_row;
    type kernel             is array ((kernel_dimension - 1) downto 0) 	    of kernel_slice_row;

end package CustomTypes;